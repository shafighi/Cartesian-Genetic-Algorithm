`timescale 1ns/1ns

module initialFsm(CLOCK_50,reset,state_controller,state_initFSM,Seed,Tap,seedIsReady,functionMemIsReady,populationCounter);//seed sefr nabashe
/*
In this function all the registers which should initial with the values of the memory will initialize.
*/
parameter population = 24;
parameter initial_controller = 2'b00;

parameter initial_initFSM = 2'b00,
			firstGenes_initFSM = 2'b01,
			popIndexSort_initFSM = 2'b10,
			finished_initFSM = 2'b11;
			
  input CLOCK_50,reset;
  input [2:0]state_controller;
  output reg [1:0]state_initFSM;
 	output reg [4095:0]Seed;
  output reg [4095:0]Tap;
	output reg seedIsReady; 
	output reg functionMemIsReady;
	output reg [7:0]populationCounter;
  //output reg initialFinished;
  
 	//initial_always
	
	

	reg start_initial,rw_initial;
  reg [19:0]address_initial;
	integer populationIndex;

  
  always@(posedge CLOCK_50)begin//initiationFSM
    if(reset)begin
		state_initFSM <= initial_initFSM;
		//initialFinished <= 0;
		Seed<=4096'd0;
		Tap<=4096'd0;
		address_initial<=20'd0;
		start_initial<=0;
		rw_initial<=0;
		seedIsReady<=0;
		functionMemIsReady<=0;
	 end else if (state_controller==initial_controller)begin 
		
			case(state_initFSM)
			
				initial_initFSM : 
				begin
					populationCounter <= 8'd0;
					Tap<=4096'h4001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
					//Seed<=4096'h5739290003040505050504784020000030100300304848400000abc0000000a7a8ac8888bbba7888800000a8000000100000001000000a658551555515550443030303005070800abbbb00000b00b0c000000d0004000404005060060060077777777777800046868056805087068706870807800000000000000000000000240486808088abbbbbbc0d00d0d0d0d0d0d0d00000ef00f0fffffffff00f0f0f0f077777777e000f000a000b00045b5b5b5b6bbbbbbbddd9d9d9f99ff7f821f1f1ff111111111111111111111111111fffffaaaaaaaaaaaaaabbbbbbbbbbbb444444444444448888888888888666666666000000003030404050696857f8f9f9f99f9f9f0f0f8f766f5f44f56666666a77a777a788888a8a888aaaaaaaaaaaaaaaaaaaaaaaaaaa653858783975874538086450386573657329876489658327573254036587325030752670828502638072654876530278028765428736528658473aaaaaaaaaaaaaaa653858783975874538086450386573657329876489658327573254036587325030752670828502638072654876530278028765428736528658473aaaaaaaaaaaaaaa653858783975874538086450386573657329876489658327573254036587325030752670828502638072654876530278028765428736528658473aaaabbbb4b4b4b4bb4b4b4bf0f0f0f0000000030003003333222fff;
					Seed<=4096'h5739290003040505050504784020000030100000304848400000abc0000000a7a8ac8088bbba7888800000a8000000100000000000000a658551555505550443030303005070800abbbb00000b00b0c000000d0004000404005060060060077777777777800046868056805087068706870807800000000000000000000000240486808088abbbbbbc0d00d0d0d0d0d0d0d00000ef00f0fffffffff00f0f0f0f077777777e000f000a000b00045b5b5b5b6bbbbbbbddd9d9d9f99ff7f821f1f1ff111111111111111111111111111fffffaaaaaaaaaaaaaabbbb1bbbbbbb441444441444448888888888888666606666000010003030404050696857f8f9f9f99f9f9f0f0f8f766f5f44f56666666a77a777a788888a8a888aaaaaaaaaaaaaaaaaaaaaaaaaaa653858783975874538086450386573657329876489658327573254036587325030752670828502638072654876530278028765428736528658473aaaaaaaaaaaaaaa653858783975874538086450386573657329876489658327573254036587325030752670828502638072654876530278028765428736528658473aaaaaaaaaaaaaaa6538587839758745380864503865736573298764896583275000000001073254036587325030752670828000000001050263807265487653027802876658473aaaabbbb4b4b4b4bb4b4b4bf0f0f0f000000003000300;
					seedIsReady <= 1;
					state_initFSM<=firstGenes_initFSM;
				end
		
				firstGenes_initFSM :
					begin
					  functionMemIsReady<=1;
					    if(population==populationCounter+1)begin
							//evalReset <= 0;
							//initialFinished <= 1; 
							 state_initFSM <= finished_initFSM;
						  end else
						   state_initFSM <= popIndexSort_initFSM;
					end
					
				popIndexSort_initFSM : 
					begin 
						populationCounter<=populationCounter+8'd1;
						state_initFSM <= firstGenes_initFSM;
					end
				finished_initFSM:
				begin
				  end
		default: 
		begin
		end					
		endcase
		end else begin //if
			//initialFinished <= 0;
			state_initFSM <= initial_initFSM;
		end
		end//always
		
	endmodule
		